// Code your testbench here
// or browse Examples
`include "uvm_macros.svh"
`include "top.sv"